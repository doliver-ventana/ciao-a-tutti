//Hello World

module HelloWorld;

  $display("Hello World");

endmodule