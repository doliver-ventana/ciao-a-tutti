//Hello World

module HelloWorld;

  //I think this is on FirstBranch
  $display("Hello World");
  //Another Comment

endmodule